//Sine wave generator
