//Top Level for Project
